package shared_pkg;
	parameter FIFO_WIDTH    = 16;
    parameter FIFO_DEPTH    = 8;
    parameter max_fifo_addr = $clog2(FIFO_DEPTH);
endpackage  